
module VerilogTest (a, b, c);

input a;
input b;
output c;
// input a, b;
// output c;

and inst1 (c, a, b);

endmodule

